-- ***********************************************************************
--
-- The ESPAM Software Tool 
-- Copyright (c) 2004-2008 Leiden University (LERC group at LIACS).
-- All rights reserved.
--
-- The use and distribution terms for this software are covered by the 
-- Common Public License 1.0 (http://opensource.org/licenses/cpl1.0.txt)
-- which can be found in the file LICENSE at the root of this distribution.
-- By using this software in any fashion, you are agreeing to be bound by 
-- the terms of this license.
--
-- You must not remove this notice, or any other, from this software.
--
-- ************************************************************************

 --
-- clocks_dcm1.vhd - clock generator module for ZBT design, using
--                   Virtex-II DCMs
--
--                   Generates 1 SSRAM clocks.
--
-- (c) Alpha Data Parallel Systems Ltd. 1999-2001
--
-- Example program for ADM-XRCIIPro-Lite
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_unsigned.all;

entity myclkrst is
    generic(
        num_clock     : integer := 2);
    port(
	    -- clocks and reset from local bus
	    lreset_l      : in    std_logic;
        lclk          : in    std_logic;
        mclk          : in    std_logic;
	    -- differential clock = 125 MHz	
	    mgt_clk       : in    std_logic;
	    mgt_clkb      : in    std_logic;
		-- control signals to the module
		ctrl          : in std_logic_vector(63 downto 0); 
		-- resets generated by the module 
		rst_power_on  : out   std_logic;
        rst_ppc1      : out   std_logic;
        rst_ppc2      : out   std_logic;
        rst_design    : out   std_logic;
		-- clocks generated by the module		
        mclk_gen      : out   std_logic;
		lclk_gen	  :	out   std_logic;
	    mgt_clk_gen   : out   std_logic;		
        clk_gen       : out   std_logic_vector(num_clock - 1 downto 0);
		-- feedback clocks
		clk_fb        : in    std_logic_vector(num_clock - 1 downto 0);
		
		locked        : out   std_logic_vector(31 downto 0));
end myclkrst;

architecture synthesis of myclkrst is

    signal sl_rst_bufg     : std_logic;
	
	signal sl_mclk_ibufg   : std_logic;
    signal sl_mclk_bufg0   : std_logic;
	signal sl_mclk_dcm0    : std_logic;
	signal sl_locked_mclk  : std_logic;
	
    signal sl_lclk_ibufg   : std_logic;
    signal sl_lclk_bufg0   : std_logic;
	signal sl_lclk_dcm0    : std_logic;
	signal sl_locked_lclk  : std_logic;	
    signal sl_rst_lclk     : std_logic;	
	
	signal sl_mgt_clk_ibufg   : std_logic;
    signal sl_mgt_clk_bufg0   : std_logic;
	signal sl_mgt_clk_dcm0    : std_logic;
	signal sl_mgt_clk_dcmfx   : std_logic;
    signal sl_mgt_clk_bufgfx  : std_logic;
	signal sl_locked_mgt_clk  : std_logic;	

	signal sl_clk_fb_ibufg  : std_logic_vector(num_clock - 1 downto 0);
    signal sl_clk_bufg0     : std_logic_vector(num_clock - 1 downto 0);
    signal sl_clk_dcm0      : std_logic_vector(num_clock - 1 downto 0);
	signal sl_locked_clk    : std_logic_vector(num_clock - 1 downto 0);
	
	signal sl_dllrst       : std_logic;
    signal sl_rstcnt       : std_logic_vector(3 downto 0);
   
    signal logic0         : std_logic;
    signal logic1         : std_logic;

    component DCM
        port(
            CLKIN         : in  std_logic;
            CLKFB         : in  std_logic;
            DSSEN         : in  std_logic;
            PSINCDEC      : in  std_logic;
            PSEN          : in  std_logic;
            PSCLK         : in  std_logic;
            RST           : in  std_logic;
            CLK0          : out std_logic;
            CLK90         : out std_logic;
            CLK180        : out std_logic;
            CLK270        : out std_logic;
            CLK2X         : out std_logic;
            CLK2X180      : out std_logic;
            CLKDV         : out std_logic;
            CLKFX         : out std_logic;
            CLKFX180      : out std_logic;
            LOCKED        : out std_logic;
            PSDONE        : out std_logic;
            STATUS        : out std_logic_vector(7 downto 0));
    end component;

    component IBUFGDS
        port (
	      O : out std_logic;
	      I : in std_logic;
	      IB: in std_logic
        );
    end component;

	component IBUFG
        port(
            I : in  std_logic;
            O : out std_logic);
    end component;
    
    component BUFG
        port(
            I : in  std_logic;
            O : out std_logic);
    end component;
	
	component FDDRRSE
	   port(
	        S : in	STD_LOGIC;
	        R : in	STD_LOGIC;
	        CE: in	STD_LOGIC;
	        D0: in	STD_LOGIC;
	        D1: in	STD_LOGIC;
	        C0: in	STD_LOGIC;
	        C1: in	STD_LOGIC;
	        Q : out	STD_LOGIC
	      );

end component;
    
    attribute DLL_FREQUENCY_MODE : string;
    attribute DUTY_CYCLE_CORRECTION : string;
    attribute STARTUP_WAIT : string;
    attribute CLK_FEEDBACK : string;
	
	attribute CLKIN_PERIOD : string;
  	attribute CLKFX_MULTIPLY : string;
  	attribute CLKFX_DIVIDE : string;
  	attribute DFS_FREQUENCY_MODE : string;

	--
    -- We can't use STARTUP_WAIT = TRUE, because we might be
    -- targetting a Virtex-II ES device.
    --
    attribute DLL_FREQUENCY_MODE of dll_lclk : label is "LOW";
    attribute DUTY_CYCLE_CORRECTION of dll_lclk : label is "TRUE";
    attribute STARTUP_WAIT of dll_lclk : label is "FALSE"; 
	
	attribute DLL_FREQUENCY_MODE of dll_mclk : label is "LOW";
    attribute DUTY_CYCLE_CORRECTION of dll_mclk : label is "TRUE";
    attribute STARTUP_WAIT of dll_mclk : label is "FALSE";	
	
	-- program dcm_mgt to produce 100MHz from 125MHz oscillator
  	attribute CLKIN_PERIOD of dll_mgt_clk   : label is "8";
  	attribute CLKFX_DIVIDE of dll_mgt_clk	: label is "5";
  	attribute CLKFX_MULTIPLY of dll_mgt_clk	: label is "4";
  	attribute DLL_FREQUENCY_MODE of dll_mgt_clk	: label is "LOW";
  	attribute DFS_FREQUENCY_MODE of dll_mgt_clk	: label is "LOW";
	
    attribute DLL_FREQUENCY_MODE of dll0 : label is "LOW";
    attribute DUTY_CYCLE_CORRECTION of dll0 : label is "TRUE";
    attribute STARTUP_WAIT of dll0 : label is "FALSE";
    attribute CLK_FEEDBACK of dll0 : label is "1X";			
	
    
begin
    
    --
    -- Define constant values
    --
    logic0 <= '0';
    logic1 <= '1';

	--
    -- Define output ports
    -- 
	
	-- all reset signals are active low ('0') 
	rst_power_on <= sl_rst_bufg;
    rst_ppc1     <= sl_rst_bufg and not ctrl(0);
    rst_ppc2     <= sl_rst_bufg and not ctrl(1);
    rst_design   <= sl_rst_bufg and not ctrl(2);
	
	mclk_gen     <= sl_mclk_bufg0;
	lclk_gen     <= sl_lclk_bufg0;
    mgt_clk_gen  <= sl_mgt_clk_bufg0;


l1:	for i in 0 to num_clock-1 generate
	  clk_gen(i) <= sl_clk_dcm0(i); 	
	end generate;	
	
	locked <= EXT(sl_locked_clk & sl_locked_mgt_clk & sl_locked_lclk & sl_locked_mclk, 32);
    
    --
    -- Use a global buffer to distribute the RESET. This avoids the
    -- problem of PAR being unable to pack registers into IOBs because
    -- various different buffered copies of the reset signal are used.
    --	
    ibufg_reset : BUFG
        port map(
            I => lreset_l,
            O => sl_rst_bufg);
			
------------------ MCLK generation module ------------------------------			
    --
    -- Input MCLK
    --
     ibufg_mclk : IBUFG
        port map(
            I => mclk,
            O => sl_mclk_ibufg); 
			    
    --
    -- Generate reset signal to DLLs/DCMs
    --
--    gen_dllrst : process(sl_rst_bufg, sl_mclk_bufg0)	  
--    begin
--        if sl_rst_bufg = '0' then
--            sl_dllrst <= '1';
--            sl_rstcnt <= (others => '0');
--        elsif sl_mclk_bufg0'event and sl_mclk_bufg0 = '1' then			
--            if sl_dllrst = '1' then
--                sl_rstcnt <= sl_rstcnt + 1;
--            end if;
--            if AND_reduce(sl_rstcnt) = '1' then
--                sl_dllrst <= '0';
--            end if;
--        end if;
--    end process;

	--
    -- Generate MCLK and derivatives
    --
    dll_mclk : DCM
        port map(
            CLKIN    => sl_mclk_ibufg,
            CLKFB    => sl_mclk_bufg0,
            DSSEN    => logic0,
            PSINCDEC => logic0,
            PSEN     => logic0,
            PSCLK    => logic0,
            RST      => logic0,
            CLK0     => sl_mclk_dcm0,
            LOCKED   => sl_locked_mclk);
		
	bufg_mclk0 : BUFG
	port map(	  
            I => sl_mclk_dcm0,
            O => sl_mclk_bufg0);
    
-------------- end MCLK generation module ------------------------------

------------------ MGT_CLK generation module ------------------------------			
    --
    -- Input MGT_CLK
    --
	ibufg_mgt_clk : IBUFGDS
	     port map (
		   I => mgt_clk,
	       IB=> mgt_clkb,
	       O => sl_mgt_clk_ibufg
    );	
	    
	--
    -- Generate MGT_CLK and derivatives
    --
    dll_mgt_clk : DCM
        port map(
            CLKIN     => sl_mgt_clk_ibufg,
            CLKFB     => sl_mgt_clk_bufg0,
            DSSEN     => logic0,
            PSINCDEC  => logic0,
            PSEN      => logic0,
            PSCLK     => logic0,
            RST       => logic0,
            CLK0      => sl_mgt_clk_dcm0,
            CLK90     => open,
            CLK180    => open,
            CLK270    => open,
            CLK2X     => open,
            CLK2X180  => open,
            CLKDV     => open,
            CLKFX     => sl_mgt_clk_dcmfx,
            CLKFX180  => open,			
            LOCKED    => sl_locked_mgt_clk, 
            PSDONE    => open,
            STATUS    => open			
			);

	bufg_mgt_clk0 : BUFG
        port map(
            I => sl_mgt_clk_dcm0,
            O => sl_mgt_clk_bufg0);
			
	bufg_mgt_clkfx : BUFG
        port map(
            I => sl_mgt_clk_dcmfx,
            O => sl_mgt_clk_bufgfx);			

-------------- end MGT_CLK generation module ------------------------------

------------------ LCLK generation module ------------------------------			
    --
    -- Input LCLK
    --
    ibufg_lclk : IBUFG
        port map(
            I => lclk,
            O => sl_lclk_ibufg);    
	--
    -- Generate LCLK and derivatives
    --
	dll_lclk : DCM
        port map(
            CLKIN    => sl_lclk_ibufg,
            CLKFB    => sl_lclk_bufg0,
            DSSEN    => logic0,
            PSINCDEC => logic0,
            PSEN     => logic0,
            PSCLK    => logic0,
            RST      => logic0,
            CLK0     => sl_lclk_dcm0,
            LOCKED   => sl_locked_lclk);
		
	bufg_lclk : BUFG
        port map(
            I => sl_lclk_dcm0,
            O => sl_lclk_bufg0);
    
-------------- end LCLK generation module ------------------------------

sl_rst_lclk <= not sl_locked_lclk;

-------------- ZBT clocks generation module ----------------------------
        
    ibufg0: IBUFG
        port map(
            I => clk_fb(0),
            O => sl_clk_fb_ibufg(0));
            
    dll0 : DCM
        port map(
            CLKIN    => sl_lclk_bufg0,
            CLKFB    => sl_clk_fb_ibufg(0),
            DSSEN    => logic0,
            PSINCDEC => logic0,
            PSEN     => logic0,
            PSCLK    => logic0,
            RST      => sl_rst_lclk,
            CLK0     => sl_clk_dcm0(0),
            LOCKED   => sl_locked_clk(0));

--fd_zbt : FDDRRSE
--   port map (
--	   S	=> '0',
--	   R	=> '0',
--	   CE	=> '1',
--	   D0	=> '1',
--	   D1	=> '0',
--	   C0	=> sl_lclk_bufg0,
--	   C1	=> not sl_lclk_bufg0,
--	   Q	=> sl_clk_dcm0(0)
--    );
			
-------------- end ZBT clocks generation module ------------------------------			

-------------- DDR clocks generation module ----------------------------------
        
    ibufg1: IBUFG
        port map(
            I => clk_fb(1),
            O => sl_clk_fb_ibufg(1));
            
    dll1 : DCM
        port map(
            CLKIN    => sl_lclk_bufg0,
            CLKFB    => sl_clk_fb_ibufg(1),
            DSSEN    => logic0,
            PSINCDEC => logic0,
            PSEN     => logic0,
            PSCLK    => logic0,
            RST      => sl_rst_lclk,
            CLK0     => sl_clk_dcm0(1),
            LOCKED   => sl_locked_clk(1));
						
-------------- end DRR clocks generation module ------------------------------	

end synthesis;
