-- ***********************************************************************
--
-- The ESPAM Software Tool 
-- Copyright (c) 2004-2008 Leiden University (LERC group at LIACS).
-- All rights reserved.
--
-- The use and distribution terms for this software are covered by the 
-- Common Public License 1.0 (http://opensource.org/licenses/cpl1.0.txt)
-- which can be found in the file LICENSE at the root of this distribution.
-- By using this software in any fashion, you are agreeing to be bound by 
-- the terms of this license.
--
-- You must not remove this notice, or any other, from this software.
--
-- ************************************************************************

-- $Id: host_design_ctrl.vhd,v 1.1 2007/12/07 22:08:31 stefanov Exp $

-- host_design_ctrl.vhd
--   Generated by wzhong

library ieee;

use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------
-- entity
-------------------------------------------------------------------------------

entity host_design_ctrl is
  generic
  (
    N_FIN  : integer                   := 1;
    PAR_WIDTH  : integer                   := 10
  );
  port
  (
    RST : in STD_LOGIC;   --RST '1' reset to 0 (stop), '0' to 1 (run);
    COMMAND_REG : in STD_LOGIC_VECTOR(31 downto 0);
    PARAMETER_REG : in STD_LOGIC_VECTOR(31 downto 0);
	FIN_REG_0 : in STD_LOGIC;
	FIN_REG_1 : in STD_LOGIC;
	FIN_REG_2 : in STD_LOGIC;
	FIN_REG_3 : in STD_LOGIC;
	FIN_REG_4 : in STD_LOGIC;
	FIN_REG_5 : in STD_LOGIC;
	FIN_REG_6 : in STD_LOGIC;
	FIN_REG_7 : in STD_LOGIC;
	FIN_REG_8 : in STD_LOGIC;
	FIN_REG_9 : in STD_LOGIC;
	FIN_REG_10 : in STD_LOGIC;
	FIN_REG_11 : in STD_LOGIC;
	FIN_REG_12 : in STD_LOGIC;
	FIN_REG_13 : in STD_LOGIC;
	FIN_REG_14 : in STD_LOGIC;
    FIN_REG_15 : in STD_LOGIC;
    FIN_REG_16 : in STD_LOGIC;
	FIN_REG_17 : in STD_LOGIC;
	FIN_REG_18 : in STD_LOGIC;
	FIN_REG_19 : in STD_LOGIC;
	RST_OUT : out STD_LOGIC;
	PARAM_DT : out STD_LOGIC_VECTOR(PAR_WIDTH-1 downto 0);
	PARAM_LD : out STD_LOGIC;
	STATUS_REG : out STD_LOGIC_VECTOR(31 downto 0)
  );
end entity host_design_ctrl;

-------------------------------------------------------------------------------
-- architecture
-------------------------------------------------------------------------------

architecture imp of host_design_ctrl is

  component host_design_ctrl_core is
    generic
    (
      N_FIN  : integer      := 1
    );
    port
    (
      RST : in STD_LOGIC;   --RST '1' reset to 0 (stop), '0' to 1 (run);
	  COMMAND_REG : in STD_LOGIC_VECTOR(31 downto 0);
	  FIN_REG : in STD_LOGIC_VECTOR(19 downto 0);
	  RST_OUT : out STD_LOGIC;
	  STATUS_REG : out STD_LOGIC_VECTOR(31 downto 0)
    );
  end component host_design_ctrl_core;

  signal sl_FIN_REG   :  std_logic_vector(19 downto 0);
-- COMMAND_REG(4) - '1' -> a parameter (from PARAMETER_REG) to be loaded into the PN

begin  ------------------------------------------------------------------------
   
   PARAM_DT <= PARAMETER_REG(PAR_WIDTH-1 downto 0);
   PARAM_LD <= COMMAND_REG(4);

  sl_FIN_REG(0) <= FIN_REG_0;
  sl_FIN_REG(1) <= FIN_REG_1;
  sl_FIN_REG(2) <= FIN_REG_2;
  sl_FIN_REG(3) <= FIN_REG_3;
  sl_FIN_REG(4) <= FIN_REG_4;
  sl_FIN_REG(5) <= FIN_REG_5;
  sl_FIN_REG(6) <= FIN_REG_6;
  sl_FIN_REG(7) <= FIN_REG_7;
  sl_FIN_REG(8) <= FIN_REG_8;
  sl_FIN_REG(9) <= FIN_REG_9;
  sl_FIN_REG(10) <= FIN_REG_10;
  sl_FIN_REG(11) <= FIN_REG_11;
  sl_FIN_REG(12) <= FIN_REG_12;
  sl_FIN_REG(13) <= FIN_REG_13;
  sl_FIN_REG(14) <= FIN_REG_14;
  sl_FIN_REG(15) <= FIN_REG_15;
  sl_FIN_REG(16) <= FIN_REG_16;
  sl_FIN_REG(17) <= FIN_REG_17;
  sl_FIN_REG(18) <= FIN_REG_18;
  sl_FIN_REG(19) <= FIN_REG_19;
	
  HOST_DESIGN_CTRL_CORE_I : host_design_ctrl_core
    generic map
    (
      N_FIN  =>  N_FIN
    )
    port map
    (
      RST           =>  RST,
      COMMAND_REG   =>  COMMAND_REG,
      FIN_REG       =>  sl_FIN_REG,
      RST_OUT       =>  RST_OUT,
      STATUS_REG    =>  STATUS_REG
    ); 

end architecture imp;

